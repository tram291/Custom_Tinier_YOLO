// system.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module system (
		input  wire        clk_50_clk,                          //     clk_50.clk
		output wire        kernel_clk_clk,                      // kernel_clk.clk
		output wire [14:0] memory_mem_a,                        //     memory.mem_a
		output wire [2:0]  memory_mem_ba,                       //           .mem_ba
		output wire        memory_mem_ck,                       //           .mem_ck
		output wire        memory_mem_ck_n,                     //           .mem_ck_n
		output wire        memory_mem_cke,                      //           .mem_cke
		output wire        memory_mem_cs_n,                     //           .mem_cs_n
		output wire        memory_mem_ras_n,                    //           .mem_ras_n
		output wire        memory_mem_cas_n,                    //           .mem_cas_n
		output wire        memory_mem_we_n,                     //           .mem_we_n
		output wire        memory_mem_reset_n,                  //           .mem_reset_n
		inout  wire [31:0] memory_mem_dq,                       //           .mem_dq
		inout  wire [3:0]  memory_mem_dqs,                      //           .mem_dqs
		inout  wire [3:0]  memory_mem_dqs_n,                    //           .mem_dqs_n
		output wire        memory_mem_odt,                      //           .mem_odt
		output wire [3:0]  memory_mem_dm,                       //           .mem_dm
		input  wire        memory_oct_rzqin,                    //           .oct_rzqin
		output wire        peripheral_hps_io_emac1_inst_TX_CLK, // peripheral.hps_io_emac1_inst_TX_CLK
		output wire        peripheral_hps_io_emac1_inst_TXD0,   //           .hps_io_emac1_inst_TXD0
		output wire        peripheral_hps_io_emac1_inst_TXD1,   //           .hps_io_emac1_inst_TXD1
		output wire        peripheral_hps_io_emac1_inst_TXD2,   //           .hps_io_emac1_inst_TXD2
		output wire        peripheral_hps_io_emac1_inst_TXD3,   //           .hps_io_emac1_inst_TXD3
		input  wire        peripheral_hps_io_emac1_inst_RXD0,   //           .hps_io_emac1_inst_RXD0
		inout  wire        peripheral_hps_io_emac1_inst_MDIO,   //           .hps_io_emac1_inst_MDIO
		output wire        peripheral_hps_io_emac1_inst_MDC,    //           .hps_io_emac1_inst_MDC
		input  wire        peripheral_hps_io_emac1_inst_RX_CTL, //           .hps_io_emac1_inst_RX_CTL
		output wire        peripheral_hps_io_emac1_inst_TX_CTL, //           .hps_io_emac1_inst_TX_CTL
		input  wire        peripheral_hps_io_emac1_inst_RX_CLK, //           .hps_io_emac1_inst_RX_CLK
		input  wire        peripheral_hps_io_emac1_inst_RXD1,   //           .hps_io_emac1_inst_RXD1
		input  wire        peripheral_hps_io_emac1_inst_RXD2,   //           .hps_io_emac1_inst_RXD2
		input  wire        peripheral_hps_io_emac1_inst_RXD3,   //           .hps_io_emac1_inst_RXD3
		inout  wire        peripheral_hps_io_sdio_inst_CMD,     //           .hps_io_sdio_inst_CMD
		inout  wire        peripheral_hps_io_sdio_inst_D0,      //           .hps_io_sdio_inst_D0
		inout  wire        peripheral_hps_io_sdio_inst_D1,      //           .hps_io_sdio_inst_D1
		output wire        peripheral_hps_io_sdio_inst_CLK,     //           .hps_io_sdio_inst_CLK
		inout  wire        peripheral_hps_io_sdio_inst_D2,      //           .hps_io_sdio_inst_D2
		inout  wire        peripheral_hps_io_sdio_inst_D3,      //           .hps_io_sdio_inst_D3
		inout  wire        peripheral_hps_io_usb1_inst_D0,      //           .hps_io_usb1_inst_D0
		inout  wire        peripheral_hps_io_usb1_inst_D1,      //           .hps_io_usb1_inst_D1
		inout  wire        peripheral_hps_io_usb1_inst_D2,      //           .hps_io_usb1_inst_D2
		inout  wire        peripheral_hps_io_usb1_inst_D3,      //           .hps_io_usb1_inst_D3
		inout  wire        peripheral_hps_io_usb1_inst_D4,      //           .hps_io_usb1_inst_D4
		inout  wire        peripheral_hps_io_usb1_inst_D5,      //           .hps_io_usb1_inst_D5
		inout  wire        peripheral_hps_io_usb1_inst_D6,      //           .hps_io_usb1_inst_D6
		inout  wire        peripheral_hps_io_usb1_inst_D7,      //           .hps_io_usb1_inst_D7
		input  wire        peripheral_hps_io_usb1_inst_CLK,     //           .hps_io_usb1_inst_CLK
		output wire        peripheral_hps_io_usb1_inst_STP,     //           .hps_io_usb1_inst_STP
		input  wire        peripheral_hps_io_usb1_inst_DIR,     //           .hps_io_usb1_inst_DIR
		input  wire        peripheral_hps_io_usb1_inst_NXT,     //           .hps_io_usb1_inst_NXT
		input  wire        peripheral_hps_io_uart0_inst_RX,     //           .hps_io_uart0_inst_RX
		output wire        peripheral_hps_io_uart0_inst_TX,     //           .hps_io_uart0_inst_TX
		inout  wire        peripheral_hps_io_i2c0_inst_SDA,     //           .hps_io_i2c0_inst_SDA
		inout  wire        peripheral_hps_io_i2c0_inst_SCL,     //           .hps_io_i2c0_inst_SCL
		inout  wire        peripheral_hps_io_gpio_inst_GPIO53,  //           .hps_io_gpio_inst_GPIO53
		input  wire        reset_50_reset_n                     //   reset_50.reset_n
	);

	wire   [63:0] avs_gemm_nn9w_cra_cra_ring_cra_master_readdata;              // gemm_ntt_jikK_system:avs_gemm_nn9W_cra_readdata -> avs_gemm_nn9W_cra_cra_ring:avm_readdata
	wire          avs_gemm_nn9w_cra_cra_ring_cra_master_read;                  // avs_gemm_nn9W_cra_cra_ring:avm_read -> gemm_ntt_jikK_system:avs_gemm_nn9W_cra_read
	wire    [4:0] avs_gemm_nn9w_cra_cra_ring_cra_master_address;               // avs_gemm_nn9W_cra_cra_ring:avm_addr -> gemm_ntt_jikK_system:avs_gemm_nn9W_cra_address
	wire    [7:0] avs_gemm_nn9w_cra_cra_ring_cra_master_byteenable;            // avs_gemm_nn9W_cra_cra_ring:avm_byteena -> gemm_ntt_jikK_system:avs_gemm_nn9W_cra_byteenable
	wire          avs_gemm_nn9w_cra_cra_ring_cra_master_readdatavalid;         // gemm_ntt_jikK_system:avs_gemm_nn9W_cra_readdatavalid -> avs_gemm_nn9W_cra_cra_ring:avm_readdatavalid
	wire          avs_gemm_nn9w_cra_cra_ring_cra_master_write;                 // avs_gemm_nn9W_cra_cra_ring:avm_write -> gemm_ntt_jikK_system:avs_gemm_nn9W_cra_write
	wire   [63:0] avs_gemm_nn9w_cra_cra_ring_cra_master_writedata;             // avs_gemm_nn9W_cra_cra_ring:avm_writedata -> gemm_ntt_jikK_system:avs_gemm_nn9W_cra_writedata
	wire   [63:0] avs_gemm_nnfw_cra_cra_ring_cra_master_readdata;              // gemm_ntt_jikK_system:avs_gemm_nnfW_cra_readdata -> avs_gemm_nnfW_cra_cra_ring:avm_readdata
	wire          avs_gemm_nnfw_cra_cra_ring_cra_master_read;                  // avs_gemm_nnfW_cra_cra_ring:avm_read -> gemm_ntt_jikK_system:avs_gemm_nnfW_cra_read
	wire    [4:0] avs_gemm_nnfw_cra_cra_ring_cra_master_address;               // avs_gemm_nnfW_cra_cra_ring:avm_addr -> gemm_ntt_jikK_system:avs_gemm_nnfW_cra_address
	wire    [7:0] avs_gemm_nnfw_cra_cra_ring_cra_master_byteenable;            // avs_gemm_nnfW_cra_cra_ring:avm_byteena -> gemm_ntt_jikK_system:avs_gemm_nnfW_cra_byteenable
	wire          avs_gemm_nnfw_cra_cra_ring_cra_master_readdatavalid;         // gemm_ntt_jikK_system:avs_gemm_nnfW_cra_readdatavalid -> avs_gemm_nnfW_cra_cra_ring:avm_readdatavalid
	wire          avs_gemm_nnfw_cra_cra_ring_cra_master_write;                 // avs_gemm_nnfW_cra_cra_ring:avm_write -> gemm_ntt_jikK_system:avs_gemm_nnfW_cra_write
	wire   [63:0] avs_gemm_nnfw_cra_cra_ring_cra_master_writedata;             // avs_gemm_nnfW_cra_cra_ring:avm_writedata -> gemm_ntt_jikK_system:avs_gemm_nnfW_cra_writedata
	wire          acl_iface_kernel_clk_clk;                                    // acl_iface:kernel_clk_clk -> [avs_gemm_nn9W_cra_cra_ring:clk, avs_gemm_nnfW_cra_cra_ring:clk, cra_root:clk, gemm_ntt_jikK_system:clock, irq_mapper:clk, mm_interconnect_0:acl_iface_kernel_clk_clk, mm_interconnect_3:acl_iface_kernel_clk_clk, rst_controller:clk]
	wire          acl_iface_kernel_clk2x_clk;                                  // acl_iface:kernel_clk2x_clk -> gemm_ntt_jikK_system:clock2x
	wire          cra_root_ring_out_datavalid;                                 // cra_root:ro_datavalid -> avs_gemm_nn9W_cra_cra_ring:ri_datavalid
	wire          cra_root_ring_out_read;                                      // cra_root:ro_read -> avs_gemm_nn9W_cra_cra_ring:ri_read
	wire   [63:0] cra_root_ring_out_data;                                      // cra_root:ro_data -> avs_gemm_nn9W_cra_cra_ring:ri_data
	wire    [5:0] cra_root_ring_out_addr;                                      // cra_root:ro_addr -> avs_gemm_nn9W_cra_cra_ring:ri_addr
	wire          cra_root_ring_out_write;                                     // cra_root:ro_write -> avs_gemm_nn9W_cra_cra_ring:ri_write
	wire    [7:0] cra_root_ring_out_byteena;                                   // cra_root:ro_byteena -> avs_gemm_nn9W_cra_cra_ring:ri_byteena
	wire          avs_gemm_nn9w_cra_cra_ring_ring_out_datavalid;               // avs_gemm_nn9W_cra_cra_ring:ro_datavalid -> avs_gemm_nnfW_cra_cra_ring:ri_datavalid
	wire          avs_gemm_nn9w_cra_cra_ring_ring_out_read;                    // avs_gemm_nn9W_cra_cra_ring:ro_read -> avs_gemm_nnfW_cra_cra_ring:ri_read
	wire   [63:0] avs_gemm_nn9w_cra_cra_ring_ring_out_data;                    // avs_gemm_nn9W_cra_cra_ring:ro_data -> avs_gemm_nnfW_cra_cra_ring:ri_data
	wire    [5:0] avs_gemm_nn9w_cra_cra_ring_ring_out_addr;                    // avs_gemm_nn9W_cra_cra_ring:ro_addr -> avs_gemm_nnfW_cra_cra_ring:ri_addr
	wire          avs_gemm_nn9w_cra_cra_ring_ring_out_write;                   // avs_gemm_nn9W_cra_cra_ring:ro_write -> avs_gemm_nnfW_cra_cra_ring:ri_write
	wire    [7:0] avs_gemm_nn9w_cra_cra_ring_ring_out_byteena;                 // avs_gemm_nn9W_cra_cra_ring:ro_byteena -> avs_gemm_nnfW_cra_cra_ring:ri_byteena
	wire          avs_gemm_nnfw_cra_cra_ring_ring_out_datavalid;               // avs_gemm_nnfW_cra_cra_ring:ro_datavalid -> cra_root:ri_datavalid
	wire          avs_gemm_nnfw_cra_cra_ring_ring_out_read;                    // avs_gemm_nnfW_cra_cra_ring:ro_read -> cra_root:ri_read
	wire   [63:0] avs_gemm_nnfw_cra_cra_ring_ring_out_data;                    // avs_gemm_nnfW_cra_cra_ring:ro_data -> cra_root:ri_data
	wire    [5:0] avs_gemm_nnfw_cra_cra_ring_ring_out_addr;                    // avs_gemm_nnfW_cra_cra_ring:ro_addr -> cra_root:ri_addr
	wire          avs_gemm_nnfw_cra_cra_ring_ring_out_write;                   // avs_gemm_nnfW_cra_cra_ring:ro_write -> cra_root:ri_write
	wire    [7:0] avs_gemm_nnfw_cra_cra_ring_ring_out_byteena;                 // avs_gemm_nnfW_cra_cra_ring:ro_byteena -> cra_root:ri_byteena
	wire          acl_iface_kernel_reset_reset;                                // acl_iface:kernel_reset_reset_n -> [avs_gemm_nn9W_cra_cra_ring:rst_n, avs_gemm_nnfW_cra_cra_ring:rst_n, cra_root:rst_n, gemm_ntt_jikK_system:resetn, mm_interconnect_0:gemm_ntt_jikK_system_clock_reset_reset_reset_bridge_in_reset_reset, mm_interconnect_3:cra_root_reset_reset_bridge_in_reset_reset]
	wire  [255:0] gemm_ntt_jikk_system_avm_memgmem0_port_0_0_rw_readdata;      // mm_interconnect_0:gemm_ntt_jikK_system_avm_memgmem0_port_0_0_rw_readdata -> gemm_ntt_jikK_system:avm_memgmem0_port_0_0_rw_readdata
	wire          gemm_ntt_jikk_system_avm_memgmem0_port_0_0_rw_waitrequest;   // mm_interconnect_0:gemm_ntt_jikK_system_avm_memgmem0_port_0_0_rw_waitrequest -> gemm_ntt_jikK_system:avm_memgmem0_port_0_0_rw_waitrequest
	wire   [29:0] gemm_ntt_jikk_system_avm_memgmem0_port_0_0_rw_address;       // gemm_ntt_jikK_system:avm_memgmem0_port_0_0_rw_address -> mm_interconnect_0:gemm_ntt_jikK_system_avm_memgmem0_port_0_0_rw_address
	wire   [31:0] gemm_ntt_jikk_system_avm_memgmem0_port_0_0_rw_byteenable;    // gemm_ntt_jikK_system:avm_memgmem0_port_0_0_rw_byteenable -> mm_interconnect_0:gemm_ntt_jikK_system_avm_memgmem0_port_0_0_rw_byteenable
	wire          gemm_ntt_jikk_system_avm_memgmem0_port_0_0_rw_read;          // gemm_ntt_jikK_system:avm_memgmem0_port_0_0_rw_read -> mm_interconnect_0:gemm_ntt_jikK_system_avm_memgmem0_port_0_0_rw_read
	wire          gemm_ntt_jikk_system_avm_memgmem0_port_0_0_rw_readdatavalid; // mm_interconnect_0:gemm_ntt_jikK_system_avm_memgmem0_port_0_0_rw_readdatavalid -> gemm_ntt_jikK_system:avm_memgmem0_port_0_0_rw_readdatavalid
	wire          gemm_ntt_jikk_system_avm_memgmem0_port_0_0_rw_write;         // gemm_ntt_jikK_system:avm_memgmem0_port_0_0_rw_write -> mm_interconnect_0:gemm_ntt_jikK_system_avm_memgmem0_port_0_0_rw_write
	wire  [255:0] gemm_ntt_jikk_system_avm_memgmem0_port_0_0_rw_writedata;     // gemm_ntt_jikK_system:avm_memgmem0_port_0_0_rw_writedata -> mm_interconnect_0:gemm_ntt_jikK_system_avm_memgmem0_port_0_0_rw_writedata
	wire    [4:0] gemm_ntt_jikk_system_avm_memgmem0_port_0_0_rw_burstcount;    // gemm_ntt_jikK_system:avm_memgmem0_port_0_0_rw_burstcount -> mm_interconnect_0:gemm_ntt_jikK_system_avm_memgmem0_port_0_0_rw_burstcount
	wire  [255:0] mm_interconnect_0_acl_iface_kernel_mem0_readdata;            // acl_iface:kernel_mem0_readdata -> mm_interconnect_0:acl_iface_kernel_mem0_readdata
	wire          mm_interconnect_0_acl_iface_kernel_mem0_waitrequest;         // acl_iface:kernel_mem0_waitrequest -> mm_interconnect_0:acl_iface_kernel_mem0_waitrequest
	wire          mm_interconnect_0_acl_iface_kernel_mem0_debugaccess;         // mm_interconnect_0:acl_iface_kernel_mem0_debugaccess -> acl_iface:kernel_mem0_debugaccess
	wire   [24:0] mm_interconnect_0_acl_iface_kernel_mem0_address;             // mm_interconnect_0:acl_iface_kernel_mem0_address -> acl_iface:kernel_mem0_address
	wire          mm_interconnect_0_acl_iface_kernel_mem0_read;                // mm_interconnect_0:acl_iface_kernel_mem0_read -> acl_iface:kernel_mem0_read
	wire   [31:0] mm_interconnect_0_acl_iface_kernel_mem0_byteenable;          // mm_interconnect_0:acl_iface_kernel_mem0_byteenable -> acl_iface:kernel_mem0_byteenable
	wire          mm_interconnect_0_acl_iface_kernel_mem0_readdatavalid;       // acl_iface:kernel_mem0_readdatavalid -> mm_interconnect_0:acl_iface_kernel_mem0_readdatavalid
	wire          mm_interconnect_0_acl_iface_kernel_mem0_write;               // mm_interconnect_0:acl_iface_kernel_mem0_write -> acl_iface:kernel_mem0_write
	wire  [255:0] mm_interconnect_0_acl_iface_kernel_mem0_writedata;           // mm_interconnect_0:acl_iface_kernel_mem0_writedata -> acl_iface:kernel_mem0_writedata
	wire    [4:0] mm_interconnect_0_acl_iface_kernel_mem0_burstcount;          // mm_interconnect_0:acl_iface_kernel_mem0_burstcount -> acl_iface:kernel_mem0_burstcount
	wire          acl_iface_kernel_cra_waitrequest;                            // mm_interconnect_3:acl_iface_kernel_cra_waitrequest -> acl_iface:kernel_cra_waitrequest
	wire   [63:0] acl_iface_kernel_cra_readdata;                               // mm_interconnect_3:acl_iface_kernel_cra_readdata -> acl_iface:kernel_cra_readdata
	wire          acl_iface_kernel_cra_debugaccess;                            // acl_iface:kernel_cra_debugaccess -> mm_interconnect_3:acl_iface_kernel_cra_debugaccess
	wire   [29:0] acl_iface_kernel_cra_address;                                // acl_iface:kernel_cra_address -> mm_interconnect_3:acl_iface_kernel_cra_address
	wire          acl_iface_kernel_cra_read;                                   // acl_iface:kernel_cra_read -> mm_interconnect_3:acl_iface_kernel_cra_read
	wire    [7:0] acl_iface_kernel_cra_byteenable;                             // acl_iface:kernel_cra_byteenable -> mm_interconnect_3:acl_iface_kernel_cra_byteenable
	wire          acl_iface_kernel_cra_readdatavalid;                          // mm_interconnect_3:acl_iface_kernel_cra_readdatavalid -> acl_iface:kernel_cra_readdatavalid
	wire   [63:0] acl_iface_kernel_cra_writedata;                              // acl_iface:kernel_cra_writedata -> mm_interconnect_3:acl_iface_kernel_cra_writedata
	wire          acl_iface_kernel_cra_write;                                  // acl_iface:kernel_cra_write -> mm_interconnect_3:acl_iface_kernel_cra_write
	wire    [0:0] acl_iface_kernel_cra_burstcount;                             // acl_iface:kernel_cra_burstcount -> mm_interconnect_3:acl_iface_kernel_cra_burstcount
	wire   [63:0] mm_interconnect_3_cra_root_cra_slave_readdata;               // cra_root:avs_readdata -> mm_interconnect_3:cra_root_cra_slave_readdata
	wire          mm_interconnect_3_cra_root_cra_slave_waitrequest;            // cra_root:avs_waitrequest -> mm_interconnect_3:cra_root_cra_slave_waitrequest
	wire    [5:0] mm_interconnect_3_cra_root_cra_slave_address;                // mm_interconnect_3:cra_root_cra_slave_address -> cra_root:avs_addr
	wire          mm_interconnect_3_cra_root_cra_slave_read;                   // mm_interconnect_3:cra_root_cra_slave_read -> cra_root:avs_read
	wire    [7:0] mm_interconnect_3_cra_root_cra_slave_byteenable;             // mm_interconnect_3:cra_root_cra_slave_byteenable -> cra_root:avs_byteena
	wire          mm_interconnect_3_cra_root_cra_slave_readdatavalid;          // cra_root:avs_readdatavalid -> mm_interconnect_3:cra_root_cra_slave_readdatavalid
	wire          mm_interconnect_3_cra_root_cra_slave_write;                  // mm_interconnect_3:cra_root_cra_slave_write -> cra_root:avs_write
	wire   [63:0] mm_interconnect_3_cra_root_cra_slave_writedata;              // mm_interconnect_3:cra_root_cra_slave_writedata -> cra_root:avs_writedata
	wire          irq_mapper_receiver0_irq;                                    // gemm_ntt_jikK_system:kernel_irq -> irq_mapper:receiver0_irq
	wire    [0:0] acl_iface_kernel_irq_irq;                                    // irq_mapper:sender_irq -> acl_iface:kernel_irq_irq
	wire          rst_controller_reset_out_reset;                              // rst_controller:reset_out -> [irq_mapper:reset, mm_interconnect_0:acl_iface_global_reset_reset_bridge_in_reset_reset, mm_interconnect_0:acl_iface_kernel_mem0_translator_reset_reset_bridge_in_reset_reset, mm_interconnect_3:acl_iface_global_reset_reset_bridge_in_reset_reset, mm_interconnect_3:acl_iface_kernel_cra_translator_reset_reset_bridge_in_reset_reset]

	system_acl_iface acl_iface (
		.acl_internal_memorg_kernel_mode         (),                                                      //       acl_internal_memorg_kernel.mode
		.acl_kernel_clk_kernel_pll_locked_export (),                                                      // acl_kernel_clk_kernel_pll_locked.export
		.config_clk_clk                          (clk_50_clk),                                            //                       config_clk.clk
		.reset_n                                 (reset_50_reset_n),                                      //                     global_reset.reset_n
		.kernel_clk_clk                          (acl_iface_kernel_clk_clk),                              //                       kernel_clk.clk
		.kernel_clk2x_clk                        (acl_iface_kernel_clk2x_clk),                            //                     kernel_clk2x.clk
		.kernel_clk_snoop_clk                    (kernel_clk_clk),                                        //                 kernel_clk_snoop.clk
		.kernel_cra_waitrequest                  (acl_iface_kernel_cra_waitrequest),                      //                       kernel_cra.waitrequest
		.kernel_cra_readdata                     (acl_iface_kernel_cra_readdata),                         //                                 .readdata
		.kernel_cra_readdatavalid                (acl_iface_kernel_cra_readdatavalid),                    //                                 .readdatavalid
		.kernel_cra_burstcount                   (acl_iface_kernel_cra_burstcount),                       //                                 .burstcount
		.kernel_cra_writedata                    (acl_iface_kernel_cra_writedata),                        //                                 .writedata
		.kernel_cra_address                      (acl_iface_kernel_cra_address),                          //                                 .address
		.kernel_cra_write                        (acl_iface_kernel_cra_write),                            //                                 .write
		.kernel_cra_read                         (acl_iface_kernel_cra_read),                             //                                 .read
		.kernel_cra_byteenable                   (acl_iface_kernel_cra_byteenable),                       //                                 .byteenable
		.kernel_cra_debugaccess                  (acl_iface_kernel_cra_debugaccess),                      //                                 .debugaccess
		.kernel_irq_irq                          (acl_iface_kernel_irq_irq),                              //                       kernel_irq.irq
		.kernel_mem0_waitrequest                 (mm_interconnect_0_acl_iface_kernel_mem0_waitrequest),   //                      kernel_mem0.waitrequest
		.kernel_mem0_readdata                    (mm_interconnect_0_acl_iface_kernel_mem0_readdata),      //                                 .readdata
		.kernel_mem0_readdatavalid               (mm_interconnect_0_acl_iface_kernel_mem0_readdatavalid), //                                 .readdatavalid
		.kernel_mem0_burstcount                  (mm_interconnect_0_acl_iface_kernel_mem0_burstcount),    //                                 .burstcount
		.kernel_mem0_writedata                   (mm_interconnect_0_acl_iface_kernel_mem0_writedata),     //                                 .writedata
		.kernel_mem0_address                     (mm_interconnect_0_acl_iface_kernel_mem0_address),       //                                 .address
		.kernel_mem0_write                       (mm_interconnect_0_acl_iface_kernel_mem0_write),         //                                 .write
		.kernel_mem0_read                        (mm_interconnect_0_acl_iface_kernel_mem0_read),          //                                 .read
		.kernel_mem0_byteenable                  (mm_interconnect_0_acl_iface_kernel_mem0_byteenable),    //                                 .byteenable
		.kernel_mem0_debugaccess                 (mm_interconnect_0_acl_iface_kernel_mem0_debugaccess),   //                                 .debugaccess
		.kernel_pll_refclk_clk                   (clk_50_clk),                                            //                kernel_pll_refclk.clk
		.kernel_reset_reset_n                    (acl_iface_kernel_reset_reset),                          //                     kernel_reset.reset_n
		.memory_mem_a                            (memory_mem_a),                                          //                           memory.mem_a
		.memory_mem_ba                           (memory_mem_ba),                                         //                                 .mem_ba
		.memory_mem_ck                           (memory_mem_ck),                                         //                                 .mem_ck
		.memory_mem_ck_n                         (memory_mem_ck_n),                                       //                                 .mem_ck_n
		.memory_mem_cke                          (memory_mem_cke),                                        //                                 .mem_cke
		.memory_mem_cs_n                         (memory_mem_cs_n),                                       //                                 .mem_cs_n
		.memory_mem_ras_n                        (memory_mem_ras_n),                                      //                                 .mem_ras_n
		.memory_mem_cas_n                        (memory_mem_cas_n),                                      //                                 .mem_cas_n
		.memory_mem_we_n                         (memory_mem_we_n),                                       //                                 .mem_we_n
		.memory_mem_reset_n                      (memory_mem_reset_n),                                    //                                 .mem_reset_n
		.memory_mem_dq                           (memory_mem_dq),                                         //                                 .mem_dq
		.memory_mem_dqs                          (memory_mem_dqs),                                        //                                 .mem_dqs
		.memory_mem_dqs_n                        (memory_mem_dqs_n),                                      //                                 .mem_dqs_n
		.memory_mem_odt                          (memory_mem_odt),                                        //                                 .mem_odt
		.memory_mem_dm                           (memory_mem_dm),                                         //                                 .mem_dm
		.memory_oct_rzqin                        (memory_oct_rzqin),                                      //                                 .oct_rzqin
		.peripheral_hps_io_emac1_inst_TX_CLK     (peripheral_hps_io_emac1_inst_TX_CLK),                   //                       peripheral.hps_io_emac1_inst_TX_CLK
		.peripheral_hps_io_emac1_inst_TXD0       (peripheral_hps_io_emac1_inst_TXD0),                     //                                 .hps_io_emac1_inst_TXD0
		.peripheral_hps_io_emac1_inst_TXD1       (peripheral_hps_io_emac1_inst_TXD1),                     //                                 .hps_io_emac1_inst_TXD1
		.peripheral_hps_io_emac1_inst_TXD2       (peripheral_hps_io_emac1_inst_TXD2),                     //                                 .hps_io_emac1_inst_TXD2
		.peripheral_hps_io_emac1_inst_TXD3       (peripheral_hps_io_emac1_inst_TXD3),                     //                                 .hps_io_emac1_inst_TXD3
		.peripheral_hps_io_emac1_inst_RXD0       (peripheral_hps_io_emac1_inst_RXD0),                     //                                 .hps_io_emac1_inst_RXD0
		.peripheral_hps_io_emac1_inst_MDIO       (peripheral_hps_io_emac1_inst_MDIO),                     //                                 .hps_io_emac1_inst_MDIO
		.peripheral_hps_io_emac1_inst_MDC        (peripheral_hps_io_emac1_inst_MDC),                      //                                 .hps_io_emac1_inst_MDC
		.peripheral_hps_io_emac1_inst_RX_CTL     (peripheral_hps_io_emac1_inst_RX_CTL),                   //                                 .hps_io_emac1_inst_RX_CTL
		.peripheral_hps_io_emac1_inst_TX_CTL     (peripheral_hps_io_emac1_inst_TX_CTL),                   //                                 .hps_io_emac1_inst_TX_CTL
		.peripheral_hps_io_emac1_inst_RX_CLK     (peripheral_hps_io_emac1_inst_RX_CLK),                   //                                 .hps_io_emac1_inst_RX_CLK
		.peripheral_hps_io_emac1_inst_RXD1       (peripheral_hps_io_emac1_inst_RXD1),                     //                                 .hps_io_emac1_inst_RXD1
		.peripheral_hps_io_emac1_inst_RXD2       (peripheral_hps_io_emac1_inst_RXD2),                     //                                 .hps_io_emac1_inst_RXD2
		.peripheral_hps_io_emac1_inst_RXD3       (peripheral_hps_io_emac1_inst_RXD3),                     //                                 .hps_io_emac1_inst_RXD3
		.peripheral_hps_io_sdio_inst_CMD         (peripheral_hps_io_sdio_inst_CMD),                       //                                 .hps_io_sdio_inst_CMD
		.peripheral_hps_io_sdio_inst_D0          (peripheral_hps_io_sdio_inst_D0),                        //                                 .hps_io_sdio_inst_D0
		.peripheral_hps_io_sdio_inst_D1          (peripheral_hps_io_sdio_inst_D1),                        //                                 .hps_io_sdio_inst_D1
		.peripheral_hps_io_sdio_inst_CLK         (peripheral_hps_io_sdio_inst_CLK),                       //                                 .hps_io_sdio_inst_CLK
		.peripheral_hps_io_sdio_inst_D2          (peripheral_hps_io_sdio_inst_D2),                        //                                 .hps_io_sdio_inst_D2
		.peripheral_hps_io_sdio_inst_D3          (peripheral_hps_io_sdio_inst_D3),                        //                                 .hps_io_sdio_inst_D3
		.peripheral_hps_io_usb1_inst_D0          (peripheral_hps_io_usb1_inst_D0),                        //                                 .hps_io_usb1_inst_D0
		.peripheral_hps_io_usb1_inst_D1          (peripheral_hps_io_usb1_inst_D1),                        //                                 .hps_io_usb1_inst_D1
		.peripheral_hps_io_usb1_inst_D2          (peripheral_hps_io_usb1_inst_D2),                        //                                 .hps_io_usb1_inst_D2
		.peripheral_hps_io_usb1_inst_D3          (peripheral_hps_io_usb1_inst_D3),                        //                                 .hps_io_usb1_inst_D3
		.peripheral_hps_io_usb1_inst_D4          (peripheral_hps_io_usb1_inst_D4),                        //                                 .hps_io_usb1_inst_D4
		.peripheral_hps_io_usb1_inst_D5          (peripheral_hps_io_usb1_inst_D5),                        //                                 .hps_io_usb1_inst_D5
		.peripheral_hps_io_usb1_inst_D6          (peripheral_hps_io_usb1_inst_D6),                        //                                 .hps_io_usb1_inst_D6
		.peripheral_hps_io_usb1_inst_D7          (peripheral_hps_io_usb1_inst_D7),                        //                                 .hps_io_usb1_inst_D7
		.peripheral_hps_io_usb1_inst_CLK         (peripheral_hps_io_usb1_inst_CLK),                       //                                 .hps_io_usb1_inst_CLK
		.peripheral_hps_io_usb1_inst_STP         (peripheral_hps_io_usb1_inst_STP),                       //                                 .hps_io_usb1_inst_STP
		.peripheral_hps_io_usb1_inst_DIR         (peripheral_hps_io_usb1_inst_DIR),                       //                                 .hps_io_usb1_inst_DIR
		.peripheral_hps_io_usb1_inst_NXT         (peripheral_hps_io_usb1_inst_NXT),                       //                                 .hps_io_usb1_inst_NXT
		.peripheral_hps_io_uart0_inst_RX         (peripheral_hps_io_uart0_inst_RX),                       //                                 .hps_io_uart0_inst_RX
		.peripheral_hps_io_uart0_inst_TX         (peripheral_hps_io_uart0_inst_TX),                       //                                 .hps_io_uart0_inst_TX
		.peripheral_hps_io_i2c0_inst_SDA         (peripheral_hps_io_i2c0_inst_SDA),                       //                                 .hps_io_i2c0_inst_SDA
		.peripheral_hps_io_i2c0_inst_SCL         (peripheral_hps_io_i2c0_inst_SCL),                       //                                 .hps_io_i2c0_inst_SCL
		.peripheral_hps_io_gpio_inst_GPIO53      (peripheral_hps_io_gpio_inst_GPIO53)                     //                                 .hps_io_gpio_inst_GPIO53
	);

	cra_ring_node #(
		.ASYNC_RESET       (1),
		.SYNCHRONIZE_RESET (0),
		.RING_ADDR_W       (5),
		.CRA_ADDR_W        (5),
		.DATA_W            (64),
		.ID_W              (1),
		.ID                (32'b00000000000000000000000000000000)
	) avs_gemm_nn9w_cra_cra_ring (
		.clk               (acl_iface_kernel_clk_clk),                            //      clock.clk
		.rst_n             (acl_iface_kernel_reset_reset),                        //      reset.reset_n
		.avm_read          (avs_gemm_nn9w_cra_cra_ring_cra_master_read),          // cra_master.read
		.avm_write         (avs_gemm_nn9w_cra_cra_ring_cra_master_write),         //           .write
		.avm_addr          (avs_gemm_nn9w_cra_cra_ring_cra_master_address),       //           .address
		.avm_byteena       (avs_gemm_nn9w_cra_cra_ring_cra_master_byteenable),    //           .byteenable
		.avm_writedata     (avs_gemm_nn9w_cra_cra_ring_cra_master_writedata),     //           .writedata
		.avm_readdata      (avs_gemm_nn9w_cra_cra_ring_cra_master_readdata),      //           .readdata
		.avm_readdatavalid (avs_gemm_nn9w_cra_cra_ring_cra_master_readdatavalid), //           .readdatavalid
		.ri_read           (cra_root_ring_out_read),                              //    ring_in.read
		.ri_write          (cra_root_ring_out_write),                             //           .write
		.ri_addr           (cra_root_ring_out_addr),                              //           .addr
		.ri_data           (cra_root_ring_out_data),                              //           .data
		.ri_byteena        (cra_root_ring_out_byteena),                           //           .byteena
		.ri_datavalid      (cra_root_ring_out_datavalid),                         //           .datavalid
		.ro_read           (avs_gemm_nn9w_cra_cra_ring_ring_out_read),            //   ring_out.read
		.ro_write          (avs_gemm_nn9w_cra_cra_ring_ring_out_write),           //           .write
		.ro_addr           (avs_gemm_nn9w_cra_cra_ring_ring_out_addr),            //           .addr
		.ro_data           (avs_gemm_nn9w_cra_cra_ring_ring_out_data),            //           .data
		.ro_byteena        (avs_gemm_nn9w_cra_cra_ring_ring_out_byteena),         //           .byteena
		.ro_datavalid      (avs_gemm_nn9w_cra_cra_ring_ring_out_datavalid)        //           .datavalid
	);

	cra_ring_node #(
		.ASYNC_RESET       (1),
		.SYNCHRONIZE_RESET (0),
		.RING_ADDR_W       (5),
		.CRA_ADDR_W        (5),
		.DATA_W            (64),
		.ID_W              (1),
		.ID                (32'b00000000000000000000000000000001)
	) avs_gemm_nnfw_cra_cra_ring (
		.clk               (acl_iface_kernel_clk_clk),                            //      clock.clk
		.rst_n             (acl_iface_kernel_reset_reset),                        //      reset.reset_n
		.avm_read          (avs_gemm_nnfw_cra_cra_ring_cra_master_read),          // cra_master.read
		.avm_write         (avs_gemm_nnfw_cra_cra_ring_cra_master_write),         //           .write
		.avm_addr          (avs_gemm_nnfw_cra_cra_ring_cra_master_address),       //           .address
		.avm_byteena       (avs_gemm_nnfw_cra_cra_ring_cra_master_byteenable),    //           .byteenable
		.avm_writedata     (avs_gemm_nnfw_cra_cra_ring_cra_master_writedata),     //           .writedata
		.avm_readdata      (avs_gemm_nnfw_cra_cra_ring_cra_master_readdata),      //           .readdata
		.avm_readdatavalid (avs_gemm_nnfw_cra_cra_ring_cra_master_readdatavalid), //           .readdatavalid
		.ri_read           (avs_gemm_nn9w_cra_cra_ring_ring_out_read),            //    ring_in.read
		.ri_write          (avs_gemm_nn9w_cra_cra_ring_ring_out_write),           //           .write
		.ri_addr           (avs_gemm_nn9w_cra_cra_ring_ring_out_addr),            //           .addr
		.ri_data           (avs_gemm_nn9w_cra_cra_ring_ring_out_data),            //           .data
		.ri_byteena        (avs_gemm_nn9w_cra_cra_ring_ring_out_byteena),         //           .byteena
		.ri_datavalid      (avs_gemm_nn9w_cra_cra_ring_ring_out_datavalid),       //           .datavalid
		.ro_read           (avs_gemm_nnfw_cra_cra_ring_ring_out_read),            //   ring_out.read
		.ro_write          (avs_gemm_nnfw_cra_cra_ring_ring_out_write),           //           .write
		.ro_addr           (avs_gemm_nnfw_cra_cra_ring_ring_out_addr),            //           .addr
		.ro_data           (avs_gemm_nnfw_cra_cra_ring_ring_out_data),            //           .data
		.ro_byteena        (avs_gemm_nnfw_cra_cra_ring_ring_out_byteena),         //           .byteena
		.ro_datavalid      (avs_gemm_nnfw_cra_cra_ring_ring_out_datavalid)        //           .datavalid
	);

	cra_ring_root #(
		.ASYNC_RESET       (1),
		.SYNCHRONIZE_RESET (0),
		.ADDR_W            (5),
		.DATA_W            (64),
		.ID_W              (1),
		.ROM_EXT_W         (0),
		.ROM_ENABLE        (0)
	) cra_root (
		.clk               (acl_iface_kernel_clk_clk),                           //     clock.clk
		.rst_n             (acl_iface_kernel_reset_reset),                       //     reset.reset_n
		.avs_write         (mm_interconnect_3_cra_root_cra_slave_write),         // cra_slave.write
		.avs_addr          (mm_interconnect_3_cra_root_cra_slave_address),       //          .address
		.avs_byteena       (mm_interconnect_3_cra_root_cra_slave_byteenable),    //          .byteenable
		.avs_writedata     (mm_interconnect_3_cra_root_cra_slave_writedata),     //          .writedata
		.avs_readdata      (mm_interconnect_3_cra_root_cra_slave_readdata),      //          .readdata
		.avs_readdatavalid (mm_interconnect_3_cra_root_cra_slave_readdatavalid), //          .readdatavalid
		.avs_waitrequest   (mm_interconnect_3_cra_root_cra_slave_waitrequest),   //          .waitrequest
		.avs_read          (mm_interconnect_3_cra_root_cra_slave_read),          //          .read
		.ri_write          (avs_gemm_nnfw_cra_cra_ring_ring_out_write),          //   ring_in.write
		.ri_addr           (avs_gemm_nnfw_cra_cra_ring_ring_out_addr),           //          .addr
		.ri_byteena        (avs_gemm_nnfw_cra_cra_ring_ring_out_byteena),        //          .byteena
		.ri_data           (avs_gemm_nnfw_cra_cra_ring_ring_out_data),           //          .data
		.ri_read           (avs_gemm_nnfw_cra_cra_ring_ring_out_read),           //          .read
		.ri_datavalid      (avs_gemm_nnfw_cra_cra_ring_ring_out_datavalid),      //          .datavalid
		.ro_read           (cra_root_ring_out_read),                             //  ring_out.read
		.ro_write          (cra_root_ring_out_write),                            //          .write
		.ro_addr           (cra_root_ring_out_addr),                             //          .addr
		.ro_data           (cra_root_ring_out_data),                             //          .data
		.ro_byteena        (cra_root_ring_out_byteena),                          //          .byteena
		.ro_datavalid      (cra_root_ring_out_datavalid)                         //          .datavalid
	);

	gemm_ntt_jikK_system gemm_ntt_jikk_system (
		.clock                                  (acl_iface_kernel_clk_clk),                                    //              clock_reset.clk
		.resetn                                 (acl_iface_kernel_reset_reset),                                //        clock_reset_reset.reset_n
		.clock2x                                (acl_iface_kernel_clk2x_clk),                                  //            clock_reset2x.clk
		.avs_gemm_nn9W_cra_read                 (avs_gemm_nn9w_cra_cra_ring_cra_master_read),                  //        avs_gemm_nn9W_cra.read
		.avs_gemm_nn9W_cra_write                (avs_gemm_nn9w_cra_cra_ring_cra_master_write),                 //                         .write
		.avs_gemm_nn9W_cra_address              (avs_gemm_nn9w_cra_cra_ring_cra_master_address),               //                         .address
		.avs_gemm_nn9W_cra_writedata            (avs_gemm_nn9w_cra_cra_ring_cra_master_writedata),             //                         .writedata
		.avs_gemm_nn9W_cra_byteenable           (avs_gemm_nn9w_cra_cra_ring_cra_master_byteenable),            //                         .byteenable
		.avs_gemm_nn9W_cra_readdata             (avs_gemm_nn9w_cra_cra_ring_cra_master_readdata),              //                         .readdata
		.avs_gemm_nn9W_cra_readdatavalid        (avs_gemm_nn9w_cra_cra_ring_cra_master_readdatavalid),         //                         .readdatavalid
		.avs_gemm_nnfW_cra_read                 (avs_gemm_nnfw_cra_cra_ring_cra_master_read),                  //        avs_gemm_nnfW_cra.read
		.avs_gemm_nnfW_cra_write                (avs_gemm_nnfw_cra_cra_ring_cra_master_write),                 //                         .write
		.avs_gemm_nnfW_cra_address              (avs_gemm_nnfw_cra_cra_ring_cra_master_address),               //                         .address
		.avs_gemm_nnfW_cra_writedata            (avs_gemm_nnfw_cra_cra_ring_cra_master_writedata),             //                         .writedata
		.avs_gemm_nnfW_cra_byteenable           (avs_gemm_nnfw_cra_cra_ring_cra_master_byteenable),            //                         .byteenable
		.avs_gemm_nnfW_cra_readdata             (avs_gemm_nnfw_cra_cra_ring_cra_master_readdata),              //                         .readdata
		.avs_gemm_nnfW_cra_readdatavalid        (avs_gemm_nnfw_cra_cra_ring_cra_master_readdatavalid),         //                         .readdatavalid
		.kernel_irq                             (irq_mapper_receiver0_irq),                                    //               kernel_irq.irq
		.avm_memgmem0_port_0_0_rw_address       (gemm_ntt_jikk_system_avm_memgmem0_port_0_0_rw_address),       // avm_memgmem0_port_0_0_rw.address
		.avm_memgmem0_port_0_0_rw_byteenable    (gemm_ntt_jikk_system_avm_memgmem0_port_0_0_rw_byteenable),    //                         .byteenable
		.avm_memgmem0_port_0_0_rw_readdatavalid (gemm_ntt_jikk_system_avm_memgmem0_port_0_0_rw_readdatavalid), //                         .readdatavalid
		.avm_memgmem0_port_0_0_rw_read          (gemm_ntt_jikk_system_avm_memgmem0_port_0_0_rw_read),          //                         .read
		.avm_memgmem0_port_0_0_rw_readdata      (gemm_ntt_jikk_system_avm_memgmem0_port_0_0_rw_readdata),      //                         .readdata
		.avm_memgmem0_port_0_0_rw_write         (gemm_ntt_jikk_system_avm_memgmem0_port_0_0_rw_write),         //                         .write
		.avm_memgmem0_port_0_0_rw_writedata     (gemm_ntt_jikk_system_avm_memgmem0_port_0_0_rw_writedata),     //                         .writedata
		.avm_memgmem0_port_0_0_rw_waitrequest   (gemm_ntt_jikk_system_avm_memgmem0_port_0_0_rw_waitrequest),   //                         .waitrequest
		.avm_memgmem0_port_0_0_rw_burstcount    (gemm_ntt_jikk_system_avm_memgmem0_port_0_0_rw_burstcount)     //                         .burstcount
	);

	system_mm_interconnect_0 mm_interconnect_0 (
		.acl_iface_kernel_clk_clk                                           (acl_iface_kernel_clk_clk),                                    //                                         acl_iface_kernel_clk.clk
		.acl_iface_global_reset_reset_bridge_in_reset_reset                 (rst_controller_reset_out_reset),                              //                 acl_iface_global_reset_reset_bridge_in_reset.reset
		.acl_iface_kernel_mem0_translator_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                              // acl_iface_kernel_mem0_translator_reset_reset_bridge_in_reset.reset
		.gemm_ntt_jikK_system_clock_reset_reset_reset_bridge_in_reset_reset (~acl_iface_kernel_reset_reset),                               // gemm_ntt_jikK_system_clock_reset_reset_reset_bridge_in_reset.reset
		.gemm_ntt_jikK_system_avm_memgmem0_port_0_0_rw_address              (gemm_ntt_jikk_system_avm_memgmem0_port_0_0_rw_address),       //                gemm_ntt_jikK_system_avm_memgmem0_port_0_0_rw.address
		.gemm_ntt_jikK_system_avm_memgmem0_port_0_0_rw_waitrequest          (gemm_ntt_jikk_system_avm_memgmem0_port_0_0_rw_waitrequest),   //                                                             .waitrequest
		.gemm_ntt_jikK_system_avm_memgmem0_port_0_0_rw_burstcount           (gemm_ntt_jikk_system_avm_memgmem0_port_0_0_rw_burstcount),    //                                                             .burstcount
		.gemm_ntt_jikK_system_avm_memgmem0_port_0_0_rw_byteenable           (gemm_ntt_jikk_system_avm_memgmem0_port_0_0_rw_byteenable),    //                                                             .byteenable
		.gemm_ntt_jikK_system_avm_memgmem0_port_0_0_rw_read                 (gemm_ntt_jikk_system_avm_memgmem0_port_0_0_rw_read),          //                                                             .read
		.gemm_ntt_jikK_system_avm_memgmem0_port_0_0_rw_readdata             (gemm_ntt_jikk_system_avm_memgmem0_port_0_0_rw_readdata),      //                                                             .readdata
		.gemm_ntt_jikK_system_avm_memgmem0_port_0_0_rw_readdatavalid        (gemm_ntt_jikk_system_avm_memgmem0_port_0_0_rw_readdatavalid), //                                                             .readdatavalid
		.gemm_ntt_jikK_system_avm_memgmem0_port_0_0_rw_write                (gemm_ntt_jikk_system_avm_memgmem0_port_0_0_rw_write),         //                                                             .write
		.gemm_ntt_jikK_system_avm_memgmem0_port_0_0_rw_writedata            (gemm_ntt_jikk_system_avm_memgmem0_port_0_0_rw_writedata),     //                                                             .writedata
		.acl_iface_kernel_mem0_address                                      (mm_interconnect_0_acl_iface_kernel_mem0_address),             //                                        acl_iface_kernel_mem0.address
		.acl_iface_kernel_mem0_write                                        (mm_interconnect_0_acl_iface_kernel_mem0_write),               //                                                             .write
		.acl_iface_kernel_mem0_read                                         (mm_interconnect_0_acl_iface_kernel_mem0_read),                //                                                             .read
		.acl_iface_kernel_mem0_readdata                                     (mm_interconnect_0_acl_iface_kernel_mem0_readdata),            //                                                             .readdata
		.acl_iface_kernel_mem0_writedata                                    (mm_interconnect_0_acl_iface_kernel_mem0_writedata),           //                                                             .writedata
		.acl_iface_kernel_mem0_burstcount                                   (mm_interconnect_0_acl_iface_kernel_mem0_burstcount),          //                                                             .burstcount
		.acl_iface_kernel_mem0_byteenable                                   (mm_interconnect_0_acl_iface_kernel_mem0_byteenable),          //                                                             .byteenable
		.acl_iface_kernel_mem0_readdatavalid                                (mm_interconnect_0_acl_iface_kernel_mem0_readdatavalid),       //                                                             .readdatavalid
		.acl_iface_kernel_mem0_waitrequest                                  (mm_interconnect_0_acl_iface_kernel_mem0_waitrequest),         //                                                             .waitrequest
		.acl_iface_kernel_mem0_debugaccess                                  (mm_interconnect_0_acl_iface_kernel_mem0_debugaccess)          //                                                             .debugaccess
	);

	system_mm_interconnect_3 mm_interconnect_3 (
		.acl_iface_kernel_clk_clk                                          (acl_iface_kernel_clk_clk),                           //                                        acl_iface_kernel_clk.clk
		.acl_iface_global_reset_reset_bridge_in_reset_reset                (rst_controller_reset_out_reset),                     //                acl_iface_global_reset_reset_bridge_in_reset.reset
		.acl_iface_kernel_cra_translator_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                     // acl_iface_kernel_cra_translator_reset_reset_bridge_in_reset.reset
		.cra_root_reset_reset_bridge_in_reset_reset                        (~acl_iface_kernel_reset_reset),                      //                        cra_root_reset_reset_bridge_in_reset.reset
		.acl_iface_kernel_cra_address                                      (acl_iface_kernel_cra_address),                       //                                        acl_iface_kernel_cra.address
		.acl_iface_kernel_cra_waitrequest                                  (acl_iface_kernel_cra_waitrequest),                   //                                                            .waitrequest
		.acl_iface_kernel_cra_burstcount                                   (acl_iface_kernel_cra_burstcount),                    //                                                            .burstcount
		.acl_iface_kernel_cra_byteenable                                   (acl_iface_kernel_cra_byteenable),                    //                                                            .byteenable
		.acl_iface_kernel_cra_read                                         (acl_iface_kernel_cra_read),                          //                                                            .read
		.acl_iface_kernel_cra_readdata                                     (acl_iface_kernel_cra_readdata),                      //                                                            .readdata
		.acl_iface_kernel_cra_readdatavalid                                (acl_iface_kernel_cra_readdatavalid),                 //                                                            .readdatavalid
		.acl_iface_kernel_cra_write                                        (acl_iface_kernel_cra_write),                         //                                                            .write
		.acl_iface_kernel_cra_writedata                                    (acl_iface_kernel_cra_writedata),                     //                                                            .writedata
		.acl_iface_kernel_cra_debugaccess                                  (acl_iface_kernel_cra_debugaccess),                   //                                                            .debugaccess
		.cra_root_cra_slave_address                                        (mm_interconnect_3_cra_root_cra_slave_address),       //                                          cra_root_cra_slave.address
		.cra_root_cra_slave_write                                          (mm_interconnect_3_cra_root_cra_slave_write),         //                                                            .write
		.cra_root_cra_slave_read                                           (mm_interconnect_3_cra_root_cra_slave_read),          //                                                            .read
		.cra_root_cra_slave_readdata                                       (mm_interconnect_3_cra_root_cra_slave_readdata),      //                                                            .readdata
		.cra_root_cra_slave_writedata                                      (mm_interconnect_3_cra_root_cra_slave_writedata),     //                                                            .writedata
		.cra_root_cra_slave_byteenable                                     (mm_interconnect_3_cra_root_cra_slave_byteenable),    //                                                            .byteenable
		.cra_root_cra_slave_readdatavalid                                  (mm_interconnect_3_cra_root_cra_slave_readdatavalid), //                                                            .readdatavalid
		.cra_root_cra_slave_waitrequest                                    (mm_interconnect_3_cra_root_cra_slave_waitrequest)    //                                                            .waitrequest
	);

	system_irq_mapper irq_mapper (
		.clk           (acl_iface_kernel_clk_clk),       //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.sender_irq    (acl_iface_kernel_irq_irq)        //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_50_reset_n),              // reset_in0.reset
		.clk            (acl_iface_kernel_clk_clk),       //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_in1      (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

endmodule
